`timescale 1ns / 1ps

module Moore_model();


endmodule
