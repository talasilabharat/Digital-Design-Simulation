`timescale 1ns / 1ps

module Univrsal_shift_register();


endmodule
